.subckt CCM1 1 2 3 4 5
Et 1 2 value={(1-v(5))*v(3,4)/v(5)}
Gd 4 3 value={(1-v(5))*i(Et)/v(5)}
.ends