.subckt CPMold control current 1 2 d
+params: L=100e-6 fs=1e5 Va=0.5 Rf=1
*

* generate d2 for CCM or DCM, see Eq.(B.31)
Ed2 d2 0 table 
+ {MIN(
+ L*fs*(v(control)-va*v(d))/Rf/(v(2)),
+ 1-v(d)
+ )} (0.01,0.01) (0.99,0.99)
*

* generate inductor current slopes, see Eqs.(B.24) and (B.26) 
Em1 m1 0 value={Rf*v(1)/L/fs}
Em2 m2 0 value={Rf*v(2)/L/fs}
*

* compute duty cycle d, see Eq.(B.32)
Eduty d 0 table 
+ {
+ 2*(v(control)*(v(d)+v(d2))
+ -v(current)-v(m2)*v(d2)*v(d2)/2)
+ /(v(m1)*v(d)+2*va*(v(d)+v(d2)))
+ } (0.01,0.01) (0.99,0.99)
*
*
.ends ; end of subcircuit CPMold