.subckt basic_diode 1 2
D1 1 2 diode
.model diode d(Is=1e-12)
.ends